
`ifndef MFP_MACRO_AHB_ROM_ADDR_WIDTH
    `define MFP_MACRO_AHB_ROM_ADDR_WIDTH 11
`endif

`ifndef MFP_MACRO_AHB_ROM_INIT_RMEMH
    `define MFP_MACRO_AHB_ROM_INIT_RMEMH ""
`endif

// SIMULATION: 16
// DE1: 10, DE0-Nano: 13, DE0-CV or Basys3: 14, Nexys 4 or DE2-115: 16, DE10-Lite: 15
`ifndef MFP_MACRO_AHB_RAM_ADDR_WIDTH
    `define MFP_MACRO_AHB_RAM_ADDR_WIDTH 10
`endif

`ifndef MFP_MACRO_AHB_RAM_INIT_RMEMH
    `define MFP_MACRO_AHB_RAM_INIT_RMEMH ""
`endif

`ifndef MFP_MACRO_CLOCK_SOURCE
    `define MFP_MACRO_CLOCK_SOURCE mfp_clock_bypass
`endif

`ifndef MFP_MACRO_CLOCK_SOURCE_MODE
    `define MFP_MACRO_CLOCK_SOURCE_MODE 50
`endif

`ifndef MFP_MACRO_CURRENT_RTL_TOOL
    `define MFP_MACRO_CURRENT_RTL_TOOL ""
`endif

`ifndef MFP_MACRO_UART_PROGAM_ENABLE
    `define MFP_MACRO_UART_PROGAM_ENABLE 0
`endif

`ifndef MFP_MACRO_UART_PROGAM_CLKFRQ
    `define MFP_MACRO_UART_PROGAM_CLKFRQ 50000000
`endif

`ifndef MFP_MACRO_UART_PROGAM_BOUDRT
    `define MFP_MACRO_UART_PROGAM_BOUDRT 115200
`endif

//`define MFP_MACRO_USE_SDRAM_MEMORY
//`define MFP_MACRO_USE_AVALON_MEMORY
//`define MFP_MACRO_USE_PMOD_ALS
//`define MFP_MACRO_USE_IRQ_EIC
//`define MFP_MACRO_USE_ADC_MAX10
//`define MFP_MACRO_USE_BUSY_MEMORY
//`define MFP_MACRO_USE_1BYTE_AHB_LOADER
//`define MFP_MACRO_DEMO_CACHE_MISSES
//`define MFP_MACRO_DEMO_PIPE_BYPASS


`define DEFAULT_WIDTH_BTN       32
`define DEFAULT_WIDTH_SW        32
`define DEFAULT_WIDTH_LEDR      32
`define DEFAULT_WIDTH_LEDG      32
`define DEFAULT_WIDTH_7SEG      32
`define DEFAULT_SDRAM_ADDR_BITS 13
`define DEFAULT_SDRAM_ROW_BITS  13
`define DEFAULT_SDRAM_COL_BITS  10
`define DEFAULT_SDRAM_DQ_BITS   16
`define DEFAULT_SDRAM_DM_BITS   2
`define DEFAULT_SDRAM_BA_BITS   2
`define DEFAULT_EJTAG_MANUFID   11'b0  //11'h02;
`define DEFAULT_EJTAG_PARTNUM   16'b0  //16'hF1;

//
// bus address decoder
//
`define MFP_RESET_RAM_ADDR_MATCH    7'h7f
`define MFP_RAM_ADDR_MATCH          3'b0
`define MFP_GPIO_ADDR_MATCH         7'h7e
`define MFP_UART_ADDR_MATCH         17'h10401
`define MFP_EIC_ADDR_MATCH          17'h10402
`define MFP_ADC_MAX10_ADDR_MATCH    17'h10403
`define MFP_ALS_ADDR_MATCH          17'h10404
